(** This module is meant as the minimal dependency of extracted code. *)
Require expr.
